module valve_control(bus_in,cold_override,bus_out);
	input cold_override;
	input[0:3] bus_in;
	output[0:1] bus_out;

endmodule
