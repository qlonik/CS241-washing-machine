module Washing-machine();
endmodule
