module valve_control(
