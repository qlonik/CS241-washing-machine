module cycle_control(bus_in,timer_done,stage_bus,output_control1,next,timer_select,valve_enable);
	input[4:0] bus_in;
	input[3:0] stage_bus;
	input timer_done;
	output[3:0] output_control1;
	output next,timer_select,valve_enable;
	
endmodule

